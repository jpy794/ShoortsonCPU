module Execute (
    output [31:0] result,
    output ready,
    input execute_type,
    input [31:0] immediate_number,
    input [63:0] register_read,
    input [31:0] forwarding
);

// ALU

// Mul/Div

endmodule