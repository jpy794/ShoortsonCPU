module Fetch1 (
    output [127:0] inst,     // 2 ways, 2 instructions each block
    input [31:0] pc
    // TODO: operation type
);

// I cache
    
endmodule