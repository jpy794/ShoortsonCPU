module CPUTop (
    input logic clk, rst_n
);



endmodule