module Fetch2 (
    output [63:0] ready_inst,
    output ready,
    input p_address_valid,
    input [31:0] p_address,
    input [127:0] inst
);

endmodule