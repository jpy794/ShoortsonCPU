module Memory1 (
    output [127:0] data_read,
    input [31:0] v_address
    // TODO: operation type
);

endmodule